*mos
********************************************************************************* 
.OPTION POST=2
.hdl "q4_mos.va"
.hdl "q4_res.va"
.model mos simple_mos
.model res resistor
*Netlist********************************************************************************

X1 3 2 0 0 mos
R 4 3 1K
Vd 4 0 DC 1.8V
Vg 2 0 PULSE(0 1.8 0 10p 10p 1n 2n)
 *********************************************************************************
.tran 10p 10n
.print V(2)
.end



